`ifndef _{:UPPERNAME:}_INTF__SV_
`define _{:UPPERNAME:}_INTF__SV_

interface {:NAME:}_intf (input clk, reset);

endinterface
`endif
